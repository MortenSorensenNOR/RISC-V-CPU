`timescale 1ns / 1ps

module module_name #(

)(
    input logic clk,
    input logic rstn
);

endmodule
