`timescale 1ns/1ps

module load_store_stage (
);

    // In here there will eventually be logic for handeling sw, sh, and sb
    // (and equivelent load instructions), but for now it will simply not do
    // much and just pass the signals to the data memeory

endmodule
