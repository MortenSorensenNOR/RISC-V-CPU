`timescale 1ns / 1ps

module cpu #(
    parameter unsigned REG_NUM = 32
)(
    input logic clk,
    input logic rstn
);


endmodule;
