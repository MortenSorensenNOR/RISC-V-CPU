`timescale 1ns/1ps

module ex_stage (
);

    // ========== ALU Controller ==========

    // ========== ALU Src A ==========

    // ========== ALU Src B ==========

    // ========== ALU ==========

endmodule
